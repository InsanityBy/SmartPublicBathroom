** Profile: "SCHEMATIC1-AF"  [ D:\PKU\SmartPublicBathroom\0_Project\1_ShowerTerminal\1_SignalInput\InfraredSensor\Stimulation\Filter&Invert-PSpiceFiles\SCHEMATIC1\AF.sim ] 

** Creating circuit file "AF.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Cadence\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "E:\Cadence\cds_spb_home\cdssetup\pspTILibDir\LMC7101A.LIB" 
.lib "E:\Cadence\cds_spb_home\cdssetup\pspTILibDir\SN74CBTLV3253.lib" 
.lib "E:\Cadence\cds_spb_home\cdssetup\pspTILibDir\lmc7101.lib" 
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 1 100
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
